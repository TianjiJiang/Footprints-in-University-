LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY SNGT IS 
	PORT(CLK : IN STD_LOGIC;
		  DOUT: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		  inCLK:OUT STD_LOGIC
		  );
END;

ARCHITECTURE DACC OF SNGT IS 
	SIGNAL DOUT_R : STD_LOGIC_VECTOR (7 DOWNTO 0);
	
	BEGIN 
	DOUT <= DOUT_R;
	PROCESS (CLK)
		BEGIN 
			IF CLK'EVENT AND CLK = '1' THEN 
				IF DOUT_R >= 98 THEN 
					DOUT_R <= "00000000";
				ELSE
					DOUT_R <= DOUT_R +1;
				END IF;
			END IF;
		inCLK <= '1';
		inCLK <= '1';
		inCLK <= '1';
		inCLK <= '0';
		inCLK <= '0';
		inCLK <= '0';
	END PROCESS;
END;